module ltc2227(
           output CLK,
           input [11: 0] D,
           input OF
       );


endmodule
